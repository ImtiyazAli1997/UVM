`include "packet.sv"
`include "sequencer.sv"
`include "driver.sv"
`include "iMonitor.sv"
`include "master_agent.sv"
`include "oMonitor.sv"
`include "slave_agent.sv"
`include "scoreboard.sv"
`include "environment.sv"
`include "test.sv"

