// Code your testbench here
// or browse Examples
`include "files.sv"


module tb;
	
	initial begin
		run_test("my_test1");
	end
endmodule